module MotionEstimator_tb();
endmodule
