`include "transaction.sv"
`include "generator.sv"
`include "ME_Interface.sv"
`include "driver.sv"
`include "environment.sv"
`include "test.sv"
