module MotionEstimator();
endmodule
